// Code your design here
// Code your design here

`define NO_SLAVES 8
`define DATA_WIDTH 32
`define ADDR_WIDTH 32

`include "apb_interconnect.sv"
`include "apb_slave.sv"
`include "apb_default_slave.sv"

// Top DUT
// This consists of APB decoder and muxing logic to connect multiple slaves to same interconnect


module apb_top_dut (input pclk,
                   input presetn,
                   input [`ADDR_WIDTH-1:0] paddr,
                   input [`DATA_WIDTH-1:0] pwdata,
                   input pwrite,
                   input penable,
                   output [`DATA_WIDTH-1:0] prdata,
                   output pready,
                   output pslverr
                   );
  
  parameter NO_SLAVES = 8;
  parameter ADDR_WIDTH = 32;
  parameter DATA_WIDTH = 32;
  
  // Intermediate signals
  
  wire [`DATA_WIDTH-1:0] s_prdata [`NO_SLAVES];  // Each slave has it's own prdata signal
  wire [`NO_SLAVES-1:0] s_pready;                // Each slave has it's own pready signal

  wire [`NO_SLAVES-1:0] psel;   // Slave select signal
  wire [`NO_SLAVES-1:0] s_pslverr;              // Slave error response generated by Default slave
  
  
  // Interconnect instantiation
  apb_interconnect DECOD_MUX (.pclk(pclk),
                              .presetn(presetn),
                              .paddr(paddr),
                              .s_pready(s_pready),
                              .s_prdata(s_prdata),
                              .s_pslverr(s_pslverr),
                              .pslverr(pslverr),
                              .psel(psel),
                              .pready(pready),
                              .prdata(prdata)
                              );
  
  
  // Slaves instantiation
  
  generate for (genvar i = 0; i < `NO_SLAVES-1; i++)
  begin : SLAVE
    
    apb_slave SLAVE_INST ( .clk(pclk),
                          .rst_n(presetn),
                          .paddr(paddr),
                          .pwrite(pwrite),
                          .psel(psel[i]),
                          .penable(penable),
                          .pwdata(pwdata),
                          .prdata(s_prdata[i]),
                          .pready(s_pready[i]),
                          .pslverr(s_pslverr[i])
                         );
  end : SLAVE
  endgenerate
  
  
  // Last slave is default slave which generates only error response
  // Default slave instantiation
  apb_default_slave SLAVE_DEF_INST ( .clk(pclk),
                             .rst_n(presetn),
                             .paddr(paddr),
                             .pwrite(pwrite),
                             .psel(psel[`NO_SLAVES-1]),
                             .penable(penable),
                             .pwdata(pwdata),
                             .prdata(s_prdata[`NO_SLAVES-1]),
                             .pready(s_pready[`NO_SLAVES-1]),
                             .pslverr(s_pslverr[`NO_SLAVES-1])
                            );
  
  
  
endmodule : apb_top_dut