
// APB interconnect
module apb_interconnect (input pclk,
                         input presetn,
                         input [`ADDR_WIDTH-1:0]  paddr,
                         input  [`NO_SLAVES-1:0] s_pready ,
                         input [`DATA_WIDTH-1:0] s_prdata [`NO_SLAVES],
                         input [`NO_SLAVES-1:0] s_pslverr,   // As of now only default slave generates slave error response
                         output reg  [`NO_SLAVES-1:0] psel,
                         output pready,
                         output [`DATA_WIDTH-1:0] prdata,
                         output reg pslverr
                        );

  parameter SLAVE_START_ADDR = 16'h00_00;
  parameter SLAVE_END_ADDR = 16'h06_FC;
  
  parameter IDLE = 0, SETUP = 1, ACCESS = 2;   // APB decoder states
  
  reg [1:0] state, nxt_state;
  
  reg [`NO_SLAVES-1:0] psel_temp;
  

  // Based on the paddr generated by Master, corresponding to psel 
  // signal is asserted to select that slave
  // These psel vector is used by apb_mux logic to properly multiplexer
  // prdata, pslverr and pready signals which are input apb master
  // Controller
  
  // Address decoder
  
  always @(posedge pclk, negedge presetn) begin
    if (~presetn) begin
      psel <= 0;
      state <= IDLE;
      //pready <= 0;
      //pslverr <=0;
    end
    else state <= nxt_state;
    
  end
  
  always @(*) begin
    case (state)
      IDLE : begin 
                psel = 0;
                nxt_state = SETUP;
             end
             
      SETUP : begin 
                if(paddr > SLAVE_END_ADDR) begin
                    psel[`NO_SLAVES-1] = 1'b1;  // Default slave is selected
                    nxt_state = ACCESS;
                end
                else if (paddr <= SLAVE_END_ADDR) begin 
                   psel = 1 << paddr[11:8]; // Otherwise based paddr bits corresponding psel signal is asserted
                    nxt_state = ACCESS;
                end
                else nxt_state = SETUP;
               end
      
      ACCESS : begin
                  if (paddr > SLAVE_END_ADDR)
                     nxt_state = IDLE; 
                  else if(s_pready[paddr[11:8]])
                     nxt_state = IDLE;
               end
    endcase
  end
  
  
  
  /*
  always @(*)
    if(paddr > SLAVE_END_ADDR)
      psel[`NO_SLAVES-1] = 1'b1;  // Default slave is selected
  else psel = 1 << paddr[11:8]; // Otherwise based paddr bits corresponding psel signal is asserted
  */
  
  // For prdata muxing
  // As prdata is latched at the end of access state, it is required keep track of 
  // psel to properly mux the data onto prdata line
  always @(posedge pclk)
    psel_temp <= psel;
  
  
  // Mux logic
  //assign pready = psel & s_pready ; // Based on psel signal, pready is selected
  
  assign pready = s_pready[$clog2(psel)];
  // Selecting prdata based on the psel signal
  assign prdata = s_prdata[$clog2(psel_temp)];
  
  // As of now only default slave generates slave error response
  assign pslverr = s_pslverr[$clog2(psel)];
  
  
endmodule : apb_interconnect
